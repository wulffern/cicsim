*cicsimgen tran

.param SEED=0

.option TEMP=27

.param vdda = 1.8

*Demo of cicsim
*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3
*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}
*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  dc {AVDD}
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
R1 VDD_1V8 VX 1k m=agauss(1,0.1,3)
R2 VX VSS 1k m=agauss(1,0.1,3)
*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save i(R1) v(VX)
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit
optran 0 0 0 100p 2n 0
tran 10p 10n 1p
write
quit
.endc
.end

